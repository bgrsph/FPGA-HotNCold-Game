----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:36:50 12/22/2017 
-- Design Name: 
-- Module Name:    Conditioner - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Conditioner is
    Port ( LuckyStrike : in  STD_LOGIC);
end Conditioner;

architecture Behavioral of Conditioner is

begin
--B�t�n �nemli ifler burada olcak. 
--if counter = 5 --> LOOSE (Assigner dan Counter � input olarak alcak)

-- if lucky 2, if signal A = 1 or signal C = 1 --> HOT // if 



end Behavioral;

